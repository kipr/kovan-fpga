`timescale 1ns / 1ps

module make_mot_linear(
	input [11:0] pwm,
	output [11:0] linearized_pwm);


	always @ (posedge clk) begin

		
			case(address) begin
			
			endcase
		
	end


endmodule
